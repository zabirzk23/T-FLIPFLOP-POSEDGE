library verilog;
use verilog.vl_types.all;
entity TFLIPFLOPPOSEDGE_vlg_vec_tst is
end TFLIPFLOPPOSEDGE_vlg_vec_tst;
